module alu(
    input enable_a,  // active low
    input [7:0] a, b,
    input [3:0] lut,
    output [7:0] q,
    output [3:0] status);



endmodule
